//Testbench for 32x1 Multiplexer using teo 8x1 Multiplexer and one 4x1 Multiplexer
module mux32x1_tb;
    reg d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,s0,s1,s2,s3,s4;
    wire out;
    
    mux32x1 mux(d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,s0,s1,s2,s3,s4,out);
    
    initial begin
        d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d20=0; d21=0; d22=0; d23=0; d24=0; d25=0; d26=0; d27=0; d28=0; d29=0; d30=0; d31=0; s0=0; s1=0; s2=0; s3=0; s4=0;
        #170 $finish;
    end
    
    initial begin
        #5  s0=0; s1=0; s2=0; s3=0; s4=0;d0=1; 
        #5  s0=0; s1=0; s2=0; s3=0; s4=1;d1=1; d0=0;
        #5  s0=0; s1=0; s2=0; s3=1; s4=0;d2=1; d1=0;
        #5  s0=0; s1=0; s2=0; s3=1; s4=1;d3=1; d2=0;
        #5  s0=0; s1=0; s2=1; s3=0; s4=0;d4=1; d3=0;
        #5  s0=0; s1=0; s2=1; s3=0; s4=1;d5=1; d4=0;
        #5  s0=0; s1=0; s2=1; s3=1; s4=0;d6=1; d5=0;
        #5  s0=0; s1=0; s2=1; s3=1; s4=1;d7=1; d6=0;
        #5  s0=0; s1=1; s2=0; s3=0; s4=0;d8=1; d7=0;
        #5  s0=0; s1=1; s2=0; s3=0; s4=1;d9=1; d8=0;
        #5  s0=0; s1=1; s2=0; s3=1; s4=0;d10=1; d9=0;
        #5  s0=0; s1=1; s2=0; s3=1; s4=1;d11=1; d10=0;
        #5  s0=0; s1=1; s2=1; s3=0; s4=0;d12=1; d11=0;
        #5  s0=0; s1=1; s2=1; s3=0; s4=1;d13=1; d12=0;
        #5  s0=0; s1=1; s2=1; s3=1; s4=0;d14=1; d13=0;
        #5  s0=0; s1=1; s2=1; s3=1; s4=1;d15=1; d14=0;
        #5  s0=1; s1=0; s2=0; s3=0; s4=0;d16=1; d15=0;
        #5  s0=1; s1=0; s2=0; s3=0; s4=1;d17=1; d16=0;
        #5  s0=1; s1=0; s2=0; s3=1; s4=0;d18=1; d17=0;
        #5  s0=1; s1=0; s2=0; s3=1; s4=1;d19=1; d18=0;
        #5  s0=1; s1=0; s2=1; s3=0; s4=0;d20=1; d19=0;
        #5  s0=1; s1=0; s2=1; s3=0; s4=1;d21=1; d20=0;
        #5  s0=1; s1=0; s2=1; s3=1; s4=0;d22=1; d21=0;
        #5  s0=1; s1=0; s2=1; s3=1; s4=1;d23=1; d22=0;
        #5  s0=1; s1=1; s2=0; s3=0; s4=0;d24=1; d23=0;
        #5  s0=1; s1=1; s2=0; s3=0; s4=1;d25=1; d24=0;
        #5  s0=1; s1=1; s2=0; s3=1; s4=0;d26=1; d25=0;
        #5  s0=1; s1=1; s2=0; s3=1; s4=1;d27=1; d26=0;
        #5  s0=1; s1=1; s2=1; s3=0; s4=0;d28=1; d27=0;
        #5  s0=1; s1=1; s2=1; s3=0; s4=1;d29=1; d28=0;
        #5  s0=1; s1=1; s2=1; s3=1; s4=0;d30=1; d29=0;
        #5  s0=1; s1=1; s2=1; s3=1; s4=1;d31=1; d30=0;
    end
    
    always @ (*)
        $monitor("At time=%t, s0=%d,s1=%d,s2=%d,s3=%d,s4=%d, d0=%d,d1=%d,d2=%d,d3=%d,d4=%d,d5=%d,d6=%d,d7=%d,d8=%d,d9=%d,d10=%d,d11=%d,d12=%d,d13=%d,d14=%d,d15=%d,d16=%d,d17=%d,d18=%d,d19=%d,d20=%d,d21=%d,d22=%d,d23=%d,d24=%d,d25=%d,d26=%d,d27=%d,d28=%d,d29=%d,d30=%d,d31=%d, out=%d",$time,s0,s1,s3,s3,s4,d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,out);
endmodule
